library verilog;
use verilog.vl_types.all;
entity FSM_RGY_LIGHT_TB is
end FSM_RGY_LIGHT_TB;
